`timescale 1 ns / 10 ps

module AvgPoolMulti_tb ();

reg clk,reset;
reg [6*28*28*16-1:0] inAvg;
wire [6*14*14*16-1:0] outAvg;

localparam PERIOD = 100;

integer i;

always
	#(PERIOD/2) clk = ~clk;
	
initial begin
    #0
    clk = 1'b0;
	  reset = 1;
    inAvg = 75264'h00000000000000000000000000000000000000000000a4afaba3aed2ae59ad01a9cba23d189818c6000000000000000000000000000000000000000000000000000000000000000000000000a469afbab211b1e42b5034f3366733042cfd266800000000000000000000000000000000000000000000000000000000000000000000a4f6af5fb13b2fdc38ee3ada3aa13a9c38c934c12d38182c0c9500000000000000000000000000000000000000000000000000009b5aa5a5afaab11c33a4392b3cb63de33e2a3d2c3c1e36f33157254c1f8c0000000000000000000000000000000000000000000000000000ac28b041b0d9333439973d8d3ff24121417140cb40103d13392732122985000000000000000000000000000000000000000000000000a4afb1afae8c35b83ac13e4b40214154425d431d423041a740303cd234bc2d4300000000000000000000000000000000000000000000a469afba21f035303b0e3e8d4073415a4274430342ff41ae414640743e32386e30d918c6000000000000000000000000000000000000a2fcade4b10d341d3a4b3ed44091413241fe427b420a418a408940694095406c3d293743258c000000000000000000000000000000009925adaeaf6532c83a813ea640b14178420e41a4413940cd405c40234034405e40933e3a394b2c3100000000000000000000000000000000a665b0ac2d48391c3e0d404b40ce410340b040173f273e0b3da53e383e4c400140683f3a3a012f9f00000000000000000000000000000000ae3428e037003d953f50405b408740563f023cd439a136df36c739453bea3fa9409d40573c41345b0000000000000000000000000000a6fcb03a34173b923ecc401d40433fe73e7d3c5938c131a50000000036143bac402140eb40e63d4f38100000000000000000000000000000ad172db038d53e1b402340673fb63d73399933662ddd2b059925aa3e36083bba405640f940f93d6838600000000000000000000000000000283233ba3b703f3f403640003de039d12fe6000000009925aaa4b1d336d03ca8409140cb407c3cd237fd000000000000000000000000000028f636e23c9f3ff340693fbc3c9a36cd00000000a469ac3cb1a621c83a193e414054405b3fb53c80373200000000000000000000000000002f9238773d7f4027406d3ec03b5d335c0000a93dafd1b2372a1e38d63d963eae3f313e9c3e2c3b0d34b80000000000000000000000000000301538973cc73fbc40213e033928a594ae9db2b8b16c32e83a7b3d453dbb3e153dd23dd43c1136af260400000000000000000000000000003026389c3d363f26401a3de838dbaf04add433e439a13c793da83e053e8b3e313e103c9538a130720000000000000000000000000000000030c038c53d093fb8401e3ea93b9639803b423cc63d6e3e883ed73ee83e5a3d8d3b49356b00000000000000000000000000000000000000003249395e3d494032412c40e13f7f3d9a3e2a3ef73f493eea3f403f0a3e223b4e3575000000000000000000000000000000000000000000002ffe39533d1540164167420c41be413740b740624075405b3fc13de33b6c36f92f05000000000000000000000000000000000000000000002d9836153bbe3f984166427a422d41b8413e40dc405e3ec13cc6391734120000000000000000000000000000000000000000000000000000279f339138203c063e8c407840ee40ee40773f343d413a08348b000000000000000000000000000000000000000000000000000000000000000026ce312437173a8d3d403e8d3ea63d343aba35902ca300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a5edb048b611b8fab967b81bb576b0d7a955000000000000000000000000000000000000000000000000000000000000000000000000a594b275b8fabc45bca5bc3db9cbb60bb143b13100000000000000000000000000000000000000000000000000000000000000000000a647b276b97abccbbd8dbe0ebe11bdecbc20b6edb10eaa5e9d1e00000000000000000000000000000000000000000000000000009ca6a909b33cb983bd1fbeffc041c097c079bf9fbe76bd16b9afb2daae3d0000000000000000000000000000000000000000000000000000ad2eb5c9baf0bd5cbfcec0b6c11dc128c147c0ecc006be36badcb0a0ac0e000000000000000000000000000000000000000000000000a5edb494ba71bd2ebf24c058c08ec12ac132c09dc04dbf2abdb1bc88b95eb37900000000000000000000000000000000000000000000a594b275b9e0bda6bf63c08bc04bc053c0b6bf76be5fc009c03abe72bce6bbd1b797a955000000000000000000000000000000000000a46ab0f1b8b1bd5bbff7c047bfb1bf87bfd6bfacbd45bcfbbfc3c067be2bbd04bca2b807ae8c000000000000000000000000000000009a82af6ab7f9bc8abf19bfa6bf03be66bd36bd61bd22b978b956bd40bf59bdcbbcb9bd29b94fb03200000000000000000000000000000000a7e0b52dbba0be94bf1dbdc3bdb1bc95bb75bc08b7e62b14ad48bb71befebe88bd3abd32bb1ab57200000000000000000000000000000000b036b970be26bf16be27bd5ebd20ba20b676b4ddabab2526a84dbab4bf04bf10bdd5bd51bba4b7bc0000000000000000000000000000a86ab5ddbcebbfcdbecbbc7bbc16b95cb521afbbac28a86a00000000ba82bf04bf4fbd7fbcf6bbadb7c00000000000000000000000000000addfb8a9be68bf6dbd14ba2bbaddb829ad1ba154a0a09cec9a82ac76bbe2bfa9bee4bcb3bc23bb15b6940000000000000000000000000000af92bafabf68beeebc16bb6cbadeb5d5a18a000000009a82aca9b61fbd9bbfe2bdd8bae1bc0aba95b6ab0000000000000000000000000000b31dbc86bf40bdbaba8cbbdab92db0f800000000a594b069b7b1bba5be75be1dbba1b8ddba1cb84fb11f0000000000000000000000000000b44ebc84beecbd1abaecbc34b98ba8c10000aa9fb479b9c2bc6dbd6dbdaebc1ab9efb978b9cbb53aa85b0000000000000000000000000000b460bc81bf01bd3abc63bcc6b991b5e6b7d1ba33bc89bd78bda6bd8bbcdfbbb3b9c0b807b392ad7598380000000000000000000000000000b45ebc81bebcbda1bddbbf2bbd6cbc53bd21bd42bd56bd29bd80bd32bb49b83fb63fb261aad1a23d00000000000000000000000000000000b3f2bc24be79be7abf0fc033bfd1be31bd89bd87be4bbe92bd84bb00b8d3b8a9b4a3a79a0000000000000000000000000000000000000000b23cbab1bd65bdddbff9c0a9c0b5c0b8c026bf6fbe7fbd85bc29b9d9b70db230ac5900000000000000000000000000000000000000000000b11cb901bc13bce7bebcc03fc01fbf5ebe90bde0bd3dbbacb680b0eab0f2a926a0ec00000000000000000000000000000000000000000000acdeb613b93fbae7bc31bd98bf2cbf64be68bc33b77fb245b129abbca5b70000000000000000000000000000000000000000000000000000a284aecfb24bb78cb9c5ba5cb9c5b7bab2f7b063b125ae2ca6600000000000000000000000000000000000000000000000000000000000000000a1d1a975a7a42c002c0c2c7e26cea99aac26a8139e820000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000098c2a4d9aacfacea9efd3029332430702965000000000000000000000000000000000000000000000000000000000000000000000000987a20862fc8365839e23bdc3c2a3b2a386c345600000000000000000000000000000000000000000000000000000000000000000000990a1e4c31d439113c2b3ec63fd93ef43d003c3238832a391d2e00000000000000000000000000000000000000000000000000008f779d251fb031fa39483c8c3f5a40cc41c241c540483d923ac135122f22000000000000000000000000000000000000000000000000000095c41e6031fc39663d3b4036421a431e437f434641e9402b3e883a9c350d00000000000000000000000000000000000000000000000098c22d0c36ab3a2b3d9d40c6429843be444344084403429c40c63ec03c6936ac00000000000000000000000000000000000000000000987a208633363a053d024073424b4353443a439a432a42d9418240293fed3ee139ec29650000000000000000000000000000000000009717227a325439ae3cce4085425e430d438942b84161413b4150414d4070404c40293c3d32ba000000000000000000000000000000008d3922bc304d38343cc4405e422b42cf42b641f540cf3fc53f10405440a6402d4064407e3d43368d0000000000000000000000000000000016a02ef038153bbd3efe416b4243421840993f343dfc3c113b593cea3e773f45408640f53e8638a600000000000000000000000000000000271034663ae93dbe409541be41af402f3dab3c2737aa319e309238643e2b3fc940ce41893f933aac00000000000000000000000000009b172f1939313cbc401341644220408e3cab37e731ef2c1f00000000382a3e37402b414341c6401f3aed0000000000000000000000000000295c358a3c293ef040e241d840cb3cda348528d927e617118d399ff037d23e29403d417c41bf3fbc397a00000000000000000000000000002ca3381a3cfd400340ca41783f1a38561bf3000000008d399ae02ab039b13e73409a416d41413df2379400000000000000000000000000002de239473e6a4043410341113da8340e00000000987aa354292436053cae400d41044127401a3c81353e0000000000000000000000000000314f3abc3eb63ff440b4406c3c672ba700009d51a0272f5c37703c1e3e904070408f3fd03d0338ca286a0000000000000000000000000000319a3aee3ec93fda405a406c3c492e52a44124fd35f73acc3d4e3efd4016406a3fce3d9d3a6e3194120f000000000000000000000000000031983aeb3ed8403a40a540873d1b39cd3a203c263e1b3f63401a406a40b040443db1393a2db41c7a0000000000000000000000000000000031ab3b083ebd4035419041bc40943f643f92400f40314064409740cb40043cc2386b2175000000000000000000000000000000000000000030a43a0c3eb640704197427f41c8414740e040e74125416240b53f643cc93905301c000000000000000000000000000000000000000000002eef38533cf14016418d427b42cc429e425741e34153407e3f283c3137e02c751b11000000000000000000000000000000000000000000002d8c370e3afa3dc3403b412541644148410540be40053d5538bc30cb201a000000000000000000000000000000000000000000000000000026cd33d239133b2e3d213ef4404140b740293dd4397e33e2209300000000000000000000000000000000000000000000000000000000000000002613315137af3a3b3b983bd9398736a831d72a2218ab00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000242a2ba530b4322b31079e90aca0aa19a03d00000000000000000000000000000000000000000000000000000000000000000000000023d72c932fb331f12cc6259429972120b0e4aa5e0000000000000000000000000000000000000000000000000000000000000000000024692c782d40306fac6aa46cadc0ab80a9a4a52fae9da224941200000000000000000000000000000000000000000000000000001a88255a2cda2d7e2d47aae4b04ead5f312835cd34e03494a5a4ae99a57e00000000000000000000000000000000000000000000000000002a552e0b31352c64af84b16ea9dc316e358c38a3374c36613019ae6eaab2000000000000000000000000000000000000000000000000242a290c2d602530ad6eb3d6b05c2b86373e337e3785372838182efca200a91b0000000000000000000000000000000000000000000023d72c9327fc30a4b125b3e8b133a9d2355a35f231a2353f35a638b6373d328016a0a03d00000000000000000000000000000000000022352a0a2b92262cae5ab0d8a0342f06346d35f63769369b3534359637e9380035fca67ca8d70000000000000000000000000000000018922a322b522cfdae3db4edb39f309d367936d13558358f36c434aa329b353b368235112574ab8c00000000000000000000000000000000243327ac29ccac91b25fb3f0308337783778354b31a22fdb32ec9d70a65c2e5c377035582fbaa46c0000000000000000000000000000000029dca6082d0fb297afd897003684388736c7341125b220672c0ab270a97821903757370233c82a880000000000000000000000000000263524500800ad2daa8ea118366136d73485311f2c5b208400000000b28ca99ea9823738364335c62c3700000000000000000000000000002002ab84aa3caff020343353373934dd2b1c9b44241a9953189229abb1a22854b0d835ab358436d52e220000000000000000000000000000a696ad9aae169f1031a9369c362f308a9dfd00000000189229482ccbacaeabbab0e4341f37da36722fa30000000000000000000000000000a9c6b06fab142dbc349d37b834db2ac20000000023d72b982f062d8db162b4dab39d35c33864362b2c940000000000000000000000000000ac38b0bea488322336c535e931841c8a000028a72d5e314c2d18af96b507b32f2ede377c36ef32769eca0000000000000000000000000000ac67b0cd1cc033b5375d381d2c5029f630b131e22fa1a85cb1a0b389b2312daf36fb37f43483282894900000000000000000000000000000ac69b0caa3a8349b36c8382032642cbe2c9aaaecae3eb37cb45cb12f313937243621326026329ebf00000000000000000000000000000000ad90b1aaacbc31fd384936062f06a892af76b308b559b47f257a35ee3777365a3221a41c0000000000000000000000000000000000000000ad36b33eb0cea110370e389930a0ab6cb331b0472d48355c3616384e369d332b24aa00000000000000000000000000000000000000000000aa7bb23cb0e7a9fe31a73450345431a2344635c536df382937bd34a1309f25229d5300000000000000000000000000000000000000000000a6feaf40b172aa9c3404353d36ae36d3372d385e37e7357b30a52c1ea22e00000000000000000000000000000000000000000000000000009f44aaecadd3b096265c33443685382637ad35bd32202deaa2e500000000000000000000000000000000000000000000000000000000000000009e7ca7f8ac29acdeaabe29ac2af02df62af021569b0a00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a8ceb131b5e9b741b5deb28cb1c2aecaa909000000000000000000000000000000000000000000000000000000000000000000000000a886b2dcb74db975ba27bb0cb899b29aa6b8b10200000000000000000000000000000000000000000000000000000000000000000000a917b2c6b640b7f9b4f1b4e5b201af832e4230fe2346a9739cd600000000000000000000000000000000000000000000000000009f8baacab320b656b5cbadd0315a38a83aa436e632ac350d32c2afb0adeb0000000000000000000000000000000000000000000000000000afa4b54fb815b597a520350e3c033dc53e8f3be8372e31c8351c2a28aa9c000000000000000000000000000000000000000000000000a8ceb25db726b68b2b68392b3d133e283e7b40223dd33b3a3710398535f22e7c00000000000000000000000000000000000000000000a886b2dcb444b3a8339c3a193e9c401b4033400f407c3f403d17374e3962382e31a6a909000000000000000000000000000000000000a72bb0ddb529b1962f2839e73db94022409f409a3eff3f6c3f8e3d2835fb37f037b234c8ae64000000000000000000000000000000009d47b04fb4f5b48f35da3b843e673f293fd2402b3ec43cbd3c8a3d543b8835c43638385d36a8940000000000000000000000000000000000a950b201b48f2f9c3a5a3e5b3f643f493dfe3cdc3b9738dc37453ba439de376637a639923871315c00000000000000000000000000000000b04eb091a0e039c63cd63efa3e593cb3396837d134da30222caf39753987398738953b0438f034670000000000000000000000000000ab2bb159a48035a53b363cec3dd33c7f388733e12dac28a000000000392f39963b2a39b63c17391e35bb0000000000000000000000000000ab5ca20034eb39c43c613d0e3b81390630f2297a232c1ef49d47aec2383339223c8d3abd3c993952371f0000000000000000000000000000263834fe38443b643c2a3c8a3926352b23d3000000009d47ae8ab4d73420392d3ca53bd43c9939ac352600000000000000000000000000002f3638323a103b0c3c043b573865305700000000a886b13cb5c0b61d37183b303d103c593c5c382030970000000000000000000000000000329c392e3a1339ae3b283aa3360029470000ad5fb45eb804b70ba1e039df3d133d773cf0398c34a62975000000000000000000000000000032f6394d39273524382f37b432beb523b6bab821b89ab81ead0f388a3cb93d4b3c673912341c2db319f6000000000000000000000000000032fe3953392634b432202c7ab2bdb95fba81b9a8b5e9340a3acb3d3a3d6f3cd6396634852d04246800000000000000000000000000000000342b3a083a1036ba360030b8aee4b520b1ea34e63b2c3d8c3e7a3e263ca238d83451295e0000000000000000000000000000000000000000346f3b823cc73c1e3a903ac43aa03af73c743da53f293f853e563c03387832ab2c880000000000000000000000000000000000000000000032d63ac73d563eb53ebe3f373f62400d405740263f533d5b3b2c367d33172b9722f4000000000000000000000000000000000000000000002ffa38af3bcc3e073f70406240a940793fa83de53c45387734c32dd5280900000000000000000000000000000000000000000000000000002809346238d23b463c4f3cfe3cce3ca13b6d38ca35143008288100000000000000000000000000000000000000000000000000000000000000002734314b369238c739c8395037b43463304829f7209800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ac1ab4d2b9a2bbd7bbccba80b89ab42cac16000000000000000000000000000000000000000000000000000000000000000000000000abb9b743bc1dbdefbecdbfafbe82bcd9ba18b5bb00000000000000000000000000000000000000000000000000000000000000000000ac58b72dbca7becfc0d9c1dcc27bc150c013bcd0b9e0ad199fd80000000000000000000000000000000000000000000000000000a26fae1ab7a4bca2bf66c180c308c392c386c249c115bf0dbd81b836b1320000000000000000000000000000000000000000000000000000b2edb9abbd66bff5c1e2c305c35ac2cec293c1a5c07dbdddbd3abae7b5ba000000000000000000000000000000000000000000000000ac1ab8cebcc7bfb2c169c280c2aac2aec0bbbfbbc047c048bd28bd3dbcffb8a200000000000000000000000000000000000000000000abb9b743bd35c017c1c9c218c1d6c19bc02fbc4ebae1bea3c029bdf1bc7dbcefb9c8ac16000000000000000000000000000000000000aa1db56bbc12bf34c16bc1d8c12cc027bdaabad3b5ceaefabbedbdeebd98bb53bc4eba4eb44300000000000000000000000000000000a081b482bb50bed0c086c0f7c070be5db689a3d43344392e39b8b0c0bc21be81bc89bd30bb6eb80f00000000000000000000000000000000ad1ab968bdb6c039c037c03cbe4db783358838c43ae53a9039cdb254bd79c040be19bdebbc08b97500000000000000000000000000000000b529bce8bfe9c052bf9cbdecb82737863a0039ef36ea321832d0ba0cbe9fc08cbeaabdacbb03b8d20000000000000000000000000000ae1dba10be9cc09bbfbcbdebb82634953a4f387c353b2eed00000000bb41beaac043bdcabd10b984b6650000000000000000000000000000b23fbc0bbf8bc021bddcbc1eb3f5355336a22f432a2127c2a081b1dfbcbdbf1dbfacbcf4bbb0b6e7b0870000000000000000000000000000b495bd17c020bf42bd76bb3cb45d341b2c5d00000000a081b1f8b9f0be1fbf8bbed8bcfab90fb1682e410000000000000000000000000000b5debd2dbf49bd8dbbbcb8b5b113339a00000000abb9b4f9baf3bdadbee1be95bd3eb999292534b134930000000000000000000000000000b500bcb5bed2bd8bbae7b949b406305f0000b095b8a7bc8bbe67bfb1bfb7be67bb80b228368236e0315d0000000000000000000000000000b4e1bca2bef8be24bcffbbe2ba2eb92ebac9bd1cbed3c015c07bc073bf5fbc02b1f537ee38fb341c22a70000000000000000000000000000b4e1bca4bf2dbfa9bf94bfdcc014c01bc008c043c0b8c127c0d3bf43ba632d68382e392835012ceb00000000000000000000000000000000b376bbd6bf1bc086c0a8c146c1a7c1f0c1ddc1b3c1bac0f4bec9b88c2bd436cc375431fe0000000000000000000000000000000000000000b028b93abcb2bfa0c0c6c1bdc2bcc344c2afc189c011bc38b3de374238d7386932b800000000000000000000000000000000000000000000a8d4b48fb947bc29bce7be03bed5bf62be5ebc12b1dd38643b243a9e382a33882bc20000000000000000000000000000000000000000000029cc2cf6a638b230b458b5d4b81cb62e2ce638fa3c0f3b80391a356c30810000000000000000000000000000000000000000000000000000260831b935553522371c39e23bfa3d103d303c31398736aa3106000000000000000000000000000000000000000000000000000000000000000025623070363339113abb3bd63b1b394136f1320a2921000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    #(PERIOD)
	  reset = 0;
    #(8*PERIOD)
    for (i = 6*14*14-1; i >=0; i = i - 1) begin
		  $displayh(outAvg[i*16+:16]);
	  end
    $stop;
end
AvgPoolMulti UUT
  (
    .clk(clk),
    .reset(reset),
    .apInput(inAvg),
    .apOutput(outAvg)
  );
endmodule

